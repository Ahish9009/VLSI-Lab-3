`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:05:33 09/29/2019 
// Design Name: 
// Module Name:    lookahead16bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lookahead16bit(
    input c_in,
    input [15:0] a,
    input [15:0] b,
    output c_out,
    output [15:0] s
    );
	 
	 wire [15:0] G, P;
	 assign G = a&b;
	 assign P = a^b;
	 assign C4 = G[3]|(P[3]&G[2])|(P[3]&P[2]&G[1])|(P[3]&P[2]&P[1]&G[0])|(P[3]&P[2]&P[1]&P[0]&c_in);
	 assign C8 = G[7]|G[6]&P[7]|G[5]&P[7]&P[6]|G[4]&P[7]&P[6]&P[5]|G[3]&P[7]&P[6]&P[5]&P[4]|G[2]&P[7]&P[6]&P[5]&P[4]&P[3]|G[1]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]|G[0]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]|P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0];
	 assign C12 = G[11]|G[10]&P[11]|G[9]&P[11]&P[10]|G[8]&P[11]&P[10]&P[9]|G[7]&P[11]&P[10]&P[9]&P[8]|G[6]&P[11]&P[10]&P[9]&P[8]&P[7]|G[5]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]|G[4]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]|G[3]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]|G[2]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]|G[1]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]|G[0]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]|P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0];
	 assign c_out = G[15]|G[14]&P[15]|G[13]&P[15]&P[14]|G[12]&P[15]&P[14]&P[13]|G[11]&P[15]&P[14]&P[13]&P[12]|G[10]&P[15]&P[14]&P[13]&P[12]&P[11]|G[9]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]|G[8]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]|G[7]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]|G[6]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]|G[5]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]|G[4]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]|G[3]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]|G[2]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]|G[1]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]|G[0]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]|P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0];
	 
	wire c_8, c_12, c_16, c_4;
	lookahead4bit A1(c_in, a[3:0], b[3:0], c_4, s[3:0]);
	lookahead4bit A2(C4, a[7:4], b[7:4], c_8, s[7:4]);
	lookahead4bit A3(C8, a[11:8], b[11:8], c_12, s[11:8]);
	lookahead4bit A4(C12, a[15:12], b[15:12], c_16, s[15:12]);


endmodule
