`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:05:33 09/29/2019 
// Design Name: 
// Module Name:    lookahead16bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lookahead16bit(
    input c_in,
    input [15:0] a,
    input [15:0] b,
    output c_out,
    output [15:0] s
    );
	 
	 wire [3:0] G0, G1, G2, G3, P0, P1, P2, P3, P4;


endmodule
